library verilog;
use verilog.vl_types.all;
entity EX_3_1_vlg_vec_tst is
end EX_3_1_vlg_vec_tst;
