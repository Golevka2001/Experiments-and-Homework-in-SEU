library verilog;
use verilog.vl_types.all;
entity EX_4_vlg_vec_tst is
end EX_4_vlg_vec_tst;
